<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-8.51883,6.19759,105.41,-49.5653</PageViewport>
<gate>
<ID>2</ID>
<type>BE_JKFF_LOW_NT</type>
<position>18.5,-22</position>
<input>
<ID>J</ID>9 </input>
<input>
<ID>K</ID>9 </input>
<output>
<ID>Q</ID>3 </output>
<input>
<ID>clock</ID>10 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3</ID>
<type>AA_LABEL</type>
<position>5.5,-27.5</position>
<gparam>LABEL_TEXT clock</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>4</ID>
<type>BE_JKFF_LOW_NT</type>
<position>36,-21.5</position>
<input>
<ID>J</ID>2 </input>
<input>
<ID>K</ID>2 </input>
<output>
<ID>Q</ID>7 </output>
<input>
<ID>clock</ID>10 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6</ID>
<type>BE_JKFF_LOW_NT</type>
<position>55.5,-21.5</position>
<input>
<ID>J</ID>1 </input>
<input>
<ID>K</ID>1 </input>
<output>
<ID>Q</ID>13 </output>
<input>
<ID>clock</ID>10 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7</ID>
<type>AA_LABEL</type>
<position>19,-21.5</position>
<gparam>LABEL_TEXT Qd</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>8</ID>
<type>BE_JKFF_LOW_NT</type>
<position>86,-22.5</position>
<input>
<ID>J</ID>8 </input>
<input>
<ID>K</ID>8 </input>
<output>
<ID>Q</ID>11 </output>
<input>
<ID>clock</ID>10 </input>
<output>
<ID>nQ</ID>4 </output>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>10</ID>
<type>AA_AND2</type>
<position>28.5,-20</position>
<input>
<ID>IN_0</ID>4 </input>
<input>
<ID>IN_1</ID>3 </input>
<output>
<ID>OUT</ID>2 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>11</ID>
<type>AA_LABEL</type>
<position>36.5,-21.5</position>
<gparam>LABEL_TEXT Qc</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>12</ID>
<type>AA_AND2</type>
<position>46.5,-19.5</position>
<input>
<ID>IN_0</ID>3 </input>
<input>
<ID>IN_1</ID>7 </input>
<output>
<ID>OUT</ID>1 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>14</ID>
<type>AA_AND2</type>
<position>66.5,-17.5</position>
<input>
<ID>IN_0</ID>11 </input>
<input>
<ID>IN_1</ID>3 </input>
<output>
<ID>OUT</ID>6 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>15</ID>
<type>AA_LABEL</type>
<position>56,-21</position>
<gparam>LABEL_TEXT Qb</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>17</ID>
<type>AA_LABEL</type>
<position>86.5,-22</position>
<gparam>LABEL_TEXT Qa</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>18</ID>
<type>AE_OR2</type>
<position>72.5,-20.5</position>
<input>
<ID>IN_0</ID>6 </input>
<input>
<ID>IN_1</ID>12 </input>
<output>
<ID>OUT</ID>8 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>20</ID>
<type>BB_CLOCK</type>
<position>11.5,-27.5</position>
<output>
<ID>CLK</ID>10 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>21</ID>
<type>AA_LABEL</type>
<position>6,-19.5</position>
<gparam>LABEL_TEXT Logic 1</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>22</ID>
<type>AA_AND3</type>
<position>65,-26</position>
<input>
<ID>IN_0</ID>3 </input>
<input>
<ID>IN_1</ID>7 </input>
<input>
<ID>IN_2</ID>13 </input>
<output>
<ID>OUT</ID>12 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>24</ID>
<type>AA_TOGGLE</type>
<position>12,-20</position>
<output>
<ID>OUT_0</ID>9 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>25</ID>
<type>AA_LABEL</type>
<position>29.5,-16.5</position>
<gparam>LABEL_TEXT Q'aQd</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>26</ID>
<type>DE_TO</type>
<position>22.5,-40.5</position>
<input>
<ID>IN_0</ID>3 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Qd</lparam></gate>
<gate>
<ID>28</ID>
<type>DE_TO</type>
<position>41.5,-40.5</position>
<input>
<ID>IN_0</ID>7 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Qc</lparam></gate>
<gate>
<ID>29</ID>
<type>AA_LABEL</type>
<position>47,-22.5</position>
<gparam>LABEL_TEXT QcQd</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>30</ID>
<type>DE_TO</type>
<position>61.5,-40.5</position>
<input>
<ID>IN_0</ID>13 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Qb</lparam></gate>
<gate>
<ID>32</ID>
<type>DE_TO</type>
<position>81.5,-41</position>
<input>
<ID>IN_0</ID>11 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Qa</lparam></gate>
<gate>
<ID>33</ID>
<type>AA_LABEL</type>
<position>67.5,-14</position>
<gparam>LABEL_TEXT QaQd</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>35</ID>
<type>AA_LABEL</type>
<position>66,-30</position>
<gparam>LABEL_TEXT QbQcQd</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>1</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>49.5,-19.5,52.5,-19.5</points>
<connection>
<GID>6</GID>
<name>J</name></connection>
<connection>
<GID>12</GID>
<name>OUT</name></connection>
<intersection>51 13</intersection></hsegment>
<vsegment>
<ID>13</ID>
<points>51,-23.5,51,-19.5</points>
<intersection>-23.5 15</intersection>
<intersection>-19.5 1</intersection></vsegment>
<hsegment>
<ID>15</ID>
<points>51,-23.5,52.5,-23.5</points>
<connection>
<GID>6</GID>
<name>K</name></connection>
<intersection>51 13</intersection></hsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>31.5,-19.5,33,-19.5</points>
<connection>
<GID>4</GID>
<name>J</name></connection>
<intersection>31.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>31.5,-23.5,31.5,-19.5</points>
<connection>
<GID>10</GID>
<name>OUT</name></connection>
<intersection>-23.5 10</intersection>
<intersection>-19.5 1</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>31.5,-23.5,33,-23.5</points>
<connection>
<GID>4</GID>
<name>K</name></connection>
<intersection>31.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>20.5,-26,40.5,-26</points>
<intersection>20.5 15</intersection>
<intersection>22.5 3</intersection>
<intersection>23 6</intersection>
<intersection>40.5 5</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>22.5,-26,22.5,-20</points>
<intersection>-26 1</intersection>
<intersection>-20 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>21.5,-20,22.5,-20</points>
<connection>
<GID>2</GID>
<name>Q</name></connection>
<intersection>22.5 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>40.5,-26,40.5,-20</points>
<intersection>-26 1</intersection>
<intersection>-20 7</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>23,-26,23,-21</points>
<intersection>-26 1</intersection>
<intersection>-21 8</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>40.5,-20,43.5,-20</points>
<intersection>40.5 5</intersection>
<intersection>43.5 9</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>23,-21,25.5,-21</points>
<connection>
<GID>10</GID>
<name>IN_1</name></connection>
<intersection>23 6</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>43.5,-20,43.5,-14.5</points>
<connection>
<GID>12</GID>
<name>IN_0</name></connection>
<intersection>-20 7</intersection>
<intersection>-14.5 10</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>43.5,-14.5,62.5,-14.5</points>
<intersection>43.5 9</intersection>
<intersection>62.5 11</intersection></hsegment>
<vsegment>
<ID>11</ID>
<points>62.5,-24,62.5,-14.5</points>
<intersection>-24 14</intersection>
<intersection>-18.5 12</intersection>
<intersection>-14.5 10</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>62.5,-18.5,63.5,-18.5</points>
<connection>
<GID>14</GID>
<name>IN_1</name></connection>
<intersection>62.5 11</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>62,-24,62.5,-24</points>
<connection>
<GID>22</GID>
<name>IN_0</name></connection>
<intersection>62.5 11</intersection></hsegment>
<vsegment>
<ID>15</ID>
<points>20.5,-40.5,20.5,-26</points>
<connection>
<GID>26</GID>
<name>IN_0</name></connection>
<intersection>-26 1</intersection></vsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>23,-8.5,90.5,-8.5</points>
<intersection>23 5</intersection>
<intersection>90.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>90.5,-24.5,90.5,-8.5</points>
<intersection>-24.5 4</intersection>
<intersection>-8.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>89,-24.5,90.5,-24.5</points>
<connection>
<GID>8</GID>
<name>nQ</name></connection>
<intersection>90.5 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>23,-19,23,-8.5</points>
<intersection>-19 6</intersection>
<intersection>-8.5 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>23,-19,25.5,-19</points>
<connection>
<GID>10</GID>
<name>IN_0</name></connection>
<intersection>23 5</intersection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>69.5,-19.5,69.5,-17.5</points>
<connection>
<GID>14</GID>
<name>OUT</name></connection>
<connection>
<GID>18</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>39.5,-12.5,60.5,-12.5</points>
<intersection>39.5 6</intersection>
<intersection>42.5 3</intersection>
<intersection>60.5 5</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>42.5,-19.5,42.5,-12.5</points>
<intersection>-19.5 4</intersection>
<intersection>-12.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>39,-19.5,42.5,-19.5</points>
<connection>
<GID>4</GID>
<name>Q</name></connection>
<intersection>42.5 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>60.5,-26,60.5,-12.5</points>
<intersection>-26 7</intersection>
<intersection>-12.5 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>39.5,-40.5,39.5,-12.5</points>
<intersection>-40.5 11</intersection>
<intersection>-20.5 9</intersection>
<intersection>-12.5 1</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>60.5,-26,62,-26</points>
<connection>
<GID>22</GID>
<name>IN_1</name></connection>
<intersection>60.5 5</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>39.5,-20.5,43.5,-20.5</points>
<connection>
<GID>12</GID>
<name>IN_1</name></connection>
<intersection>39.5 6</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>39.5,-40.5,39.5,-40.5</points>
<connection>
<GID>28</GID>
<name>IN_0</name></connection>
<intersection>39.5 6</intersection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>82,-24.5,82,-20.5</points>
<intersection>-24.5 3</intersection>
<intersection>-20.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>75.5,-20.5,83,-20.5</points>
<connection>
<GID>8</GID>
<name>J</name></connection>
<connection>
<GID>18</GID>
<name>OUT</name></connection>
<intersection>82 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>82,-24.5,83,-24.5</points>
<connection>
<GID>8</GID>
<name>K</name></connection>
<intersection>82 0</intersection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>15,-24,15,-18</points>
<intersection>-24 1</intersection>
<intersection>-18 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>15,-24,15.5,-24</points>
<connection>
<GID>2</GID>
<name>K</name></connection>
<intersection>15 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>14,-18,15.5,-18</points>
<intersection>14 5</intersection>
<intersection>15 0</intersection>
<intersection>15.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>15.5,-20,15.5,-18</points>
<intersection>-20 8</intersection>
<intersection>-18 2</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>14,-20,14,-18</points>
<intersection>-20 9</intersection>
<intersection>-18 2</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>15.5,-20,15.5,-20</points>
<connection>
<GID>2</GID>
<name>J</name></connection>
<intersection>15.5 4</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>14,-20,14,-20</points>
<connection>
<GID>24</GID>
<name>OUT_0</name></connection>
<intersection>14 5</intersection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>15.5,-32,83,-32</points>
<intersection>15.5 3</intersection>
<intersection>33 7</intersection>
<intersection>52.5 6</intersection>
<intersection>83 9</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>15.5,-32,15.5,-22</points>
<connection>
<GID>20</GID>
<name>CLK</name></connection>
<intersection>-32 1</intersection>
<intersection>-22 10</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>52.5,-32,52.5,-21.5</points>
<connection>
<GID>6</GID>
<name>clock</name></connection>
<intersection>-32 1</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>33,-32,33,-21.5</points>
<connection>
<GID>4</GID>
<name>clock</name></connection>
<intersection>-32 1</intersection></vsegment>
<vsegment>
<ID>9</ID>
<points>83,-32,83,-22.5</points>
<connection>
<GID>8</GID>
<name>clock</name></connection>
<intersection>-32 1</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>15.5,-22,15.5,-22</points>
<connection>
<GID>2</GID>
<name>clock</name></connection>
<intersection>15.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>63,-12,89,-12</points>
<intersection>63 3</intersection>
<intersection>89 4</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>63,-16.5,63,-12</points>
<intersection>-16.5 5</intersection>
<intersection>-12 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>89,-38,89,-12</points>
<connection>
<GID>8</GID>
<name>Q</name></connection>
<intersection>-38 6</intersection>
<intersection>-12 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>63,-16.5,63.5,-16.5</points>
<connection>
<GID>14</GID>
<name>IN_0</name></connection>
<intersection>63 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>79.5,-38,89,-38</points>
<intersection>79.5 7</intersection>
<intersection>89 4</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>79.5,-41,79.5,-38</points>
<intersection>-41 9</intersection>
<intersection>-38 6</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>79.5,-41,79.5,-41</points>
<connection>
<GID>32</GID>
<name>IN_0</name></connection>
<intersection>79.5 7</intersection></hsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>68.5,-26,68.5,-21.5</points>
<intersection>-26 1</intersection>
<intersection>-21.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>68,-26,68.5,-26</points>
<connection>
<GID>22</GID>
<name>OUT</name></connection>
<intersection>68.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>68.5,-21.5,69.5,-21.5</points>
<connection>
<GID>18</GID>
<name>IN_1</name></connection>
<intersection>68.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>59,-40.5,59,-19.5</points>
<intersection>-40.5 3</intersection>
<intersection>-28 1</intersection>
<intersection>-19.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>59,-28,62,-28</points>
<connection>
<GID>22</GID>
<name>IN_2</name></connection>
<intersection>59 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>58.5,-19.5,59,-19.5</points>
<connection>
<GID>6</GID>
<name>Q</name></connection>
<intersection>59 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>59,-40.5,59.5,-40.5</points>
<connection>
<GID>30</GID>
<name>IN_0</name></connection>
<intersection>59 0</intersection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>0,31.4959,292.996,-111.913</PageViewport></page 1>
<page 2>
<PageViewport>0,31.4959,292.996,-111.913</PageViewport></page 2>
<page 3>
<PageViewport>0,31.4959,292.996,-111.913</PageViewport></page 3>
<page 4>
<PageViewport>0,31.4959,292.996,-111.913</PageViewport></page 4>
<page 5>
<PageViewport>0,31.4959,292.996,-111.913</PageViewport></page 5>
<page 6>
<PageViewport>0,31.4959,292.996,-111.913</PageViewport></page 6>
<page 7>
<PageViewport>0,31.4959,292.996,-111.913</PageViewport></page 7>
<page 8>
<PageViewport>0,31.4959,292.996,-111.913</PageViewport></page 8>
<page 9>
<PageViewport>0,31.4959,292.996,-111.913</PageViewport></page 9></circuit>